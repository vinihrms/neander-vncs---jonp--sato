--Jump Negative