--Jump Zero