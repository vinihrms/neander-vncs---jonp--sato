--Jump