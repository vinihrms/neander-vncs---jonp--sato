--Not